*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'penatb' on Sun Feb 24 2019 at 19:01:58

*
* Globals.
*
.global GROUND VDD

*
* MAIN CELL: Component pathname : $LAB_1/Tutorials/Tutorial_5
*
        M4 Y A GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M3 Y B GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M2 Y A N$5 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M1 N$5 B VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
*
.end
