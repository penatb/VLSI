* Component: $LAB_1/Tutorials/Tutorial_5  Viewpoint: default
.INCLUDE $LAB_1/Tutorials/Tutorial_5/default/Tutorial_5_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(A)
.PROBE TRAN V(B)
.PROBE TRAN V(Y)

* --- Params
.TEMP 27
.PARAM t_sweep=0 
.STEP PARAM t_sweep 0n 100n INCR 1n

* --- Forces
VFORCE_IN A GROUND PULSE (0 2.5V 50n 1n 1n 50n 100n)
VFORCE_IN_1 B GROUND PULSE (0 2.5V 25n 1n 1n 25n 50n)
VFORCE_VDD VDD GROUND dc 2.5V

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

