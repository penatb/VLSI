*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'penatb' on Fri Feb  8 2019 at 10:41:46

*
* Globals.
*
.global GROUND VDD

*
* MAIN CELL: Component pathname : $LAB_1/Tutorials/Tutorial_1
*
        C1 OUT GROUND 2P
        M2 OUT IN VDD VDD pmos w=1.45u l=0.13u m=1 as=0.493p ad=0.493p ps=2.13u
+  pd=2.13u
        M1 OUT IN GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
*
.end
