* Component: $LAB_1/Tutorials/Tutorial_1  Viewpoint: default
.INCLUDE $LAB_1/Tutorials/Tutorial_1/default/Tutorial_1_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 200N

* --- Waveform Outputs
.PROBE TRAN V(IN)
.PROBE TRAN V(OUT)

* --- Params
.TEMP 27
.PARAM t_sweep=0 
.STEP PARAM t_sweep 0n 200n INCR 1n

* --- Forces
VFORCE__IN VDD GROUND dc 2.5V
VtsweepFORCE_IN IN GROUND PULSE (0 2.5v 25n 1n 1n 75n 150n)

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

