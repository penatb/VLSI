* Component: $LAB_1/Tutorials/Tutorial_6  Viewpoint: default
.INCLUDE $LAB_1/Tutorials/Tutorial_6/default/Tutorial_6_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(OUT)
.PROBE TRAN V(IN1)
.PROBE TRAN V(IN2)

* --- Params
.TEMP 27
.PARAM t_sweep=0 
.STEP PARAM t_sweep 0n 100n INCR 1n

* --- Forces
VFORCE__IN1 IN1 GROUND PULSE (0 2.5V 50ns 1n 1n 50n 100n)
VFORCE__IN1_1 IN2 GROUND PULSE (0 2.5V 25n 1n 1n 25n 50n)

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

